library verilog;
use verilog.vl_types.all;
entity divisiontb is
end divisiontb;

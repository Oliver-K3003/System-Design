library verilog;
use verilog.vl_types.all;
entity bidirectionalBustb is
end bidirectionalBustb;

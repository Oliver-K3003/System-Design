library verilog;
use verilog.vl_types.all;
entity multipliertb is
end multipliertb;

library verilog;
use verilog.vl_types.all;
entity control_unittb is
end control_unittb;

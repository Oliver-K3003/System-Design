`timescale 1ns/10ps

module busMUXtb;
	
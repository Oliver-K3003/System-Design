library verilog;
use verilog.vl_types.all;
entity datapath is
    port(
        HIin            : out    vl_logic;
        LOin            : out    vl_logic;
        PCin            : out    vl_logic;
        MDRin           : out    vl_logic;
        Zin             : out    vl_logic;
        Yin             : out    vl_logic;
        MARin           : out    vl_logic;
        IRin            : out    vl_logic;
        CONin           : out    vl_logic;
        OUTPORTin       : out    vl_logic;
        HIout           : out    vl_logic;
        LOout           : out    vl_logic;
        ZHIout          : out    vl_logic;
        ZLOout          : out    vl_logic;
        PCout           : out    vl_logic;
        MDRout          : out    vl_logic;
        INPORTout       : out    vl_logic;
        OUTPORTout      : out    vl_logic;
        Cout            : out    vl_logic;
        Yout            : out    vl_logic;
        Gra             : out    vl_logic;
        Grb             : out    vl_logic;
        Grc             : out    vl_logic;
        Rin             : out    vl_logic;
        Rout            : out    vl_logic;
        BAout           : out    vl_logic;
        Read            : out    vl_logic;
        IncPC           : out    vl_logic;
        write           : out    vl_logic;
        run             : out    vl_logic;
        Clock           : in     vl_logic;
        Reset           : in     vl_logic;
        Stop            : in     vl_logic;
        inportInput     : in     vl_logic_vector(31 downto 0);
        regIn           : out    vl_logic_vector(15 downto 0);
        busMuxOut       : out    vl_logic_vector(31 downto 0);
        encoderOut      : out    vl_logic_vector(4 downto 0);
        CON             : out    vl_logic;
        BusMuxInR0      : out    vl_logic_vector(31 downto 0);
        BusMuxInR1      : out    vl_logic_vector(31 downto 0);
        BusMuxInR2      : out    vl_logic_vector(31 downto 0);
        BusMuxInR3      : out    vl_logic_vector(31 downto 0);
        BusMuxInR4      : out    vl_logic_vector(31 downto 0);
        BusMuxInR5      : out    vl_logic_vector(31 downto 0);
        BusMuxInR6      : out    vl_logic_vector(31 downto 0);
        BusMuxInR7      : out    vl_logic_vector(31 downto 0);
        BusMuxInR8      : out    vl_logic_vector(31 downto 0);
        BusMuxInR9      : out    vl_logic_vector(31 downto 0);
        BusMuxInR10     : out    vl_logic_vector(31 downto 0);
        BusMuxInR11     : out    vl_logic_vector(31 downto 0);
        BusMuxInR12     : out    vl_logic_vector(31 downto 0);
        BusMuxInR13     : out    vl_logic_vector(31 downto 0);
        BusMuxInR14     : out    vl_logic_vector(31 downto 0);
        BusMuxInR15     : out    vl_logic_vector(31 downto 0);
        BusMuxInHI      : out    vl_logic_vector(31 downto 0);
        BusMuxInLO      : out    vl_logic_vector(31 downto 0);
        BusMuxInZhi     : out    vl_logic_vector(31 downto 0);
        BusMuxInZlo     : out    vl_logic_vector(31 downto 0);
        BusMuxInPC      : out    vl_logic_vector(31 downto 0);
        BusMuxInMDR     : out    vl_logic_vector(31 downto 0);
        BusMuxInInport  : out    vl_logic_vector(31 downto 0);
        BusMuxInOutport : out    vl_logic_vector(31 downto 0);
        BusMuxInY       : out    vl_logic_vector(31 downto 0);
        IRregister      : out    vl_logic_vector(31 downto 0);
        Cregister       : out    vl_logic_vector(31 downto 0);
        marToRam        : out    vl_logic_vector(8 downto 0);
        mdrToRam        : out    vl_logic_vector(31 downto 0)
    );
end datapath;

library verilog;
use verilog.vl_types.all;
entity control_unit is
    generic(
        reset_state     : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        fetch0          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        fetch1          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        fetch2          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1);
        add3            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        add4            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1);
        add5            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        sub3            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1);
        sub4            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        sub5            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1);
        mul3            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        mul4            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1);
        mul5            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0);
        mul6            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1);
        div3            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0);
        div4            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1);
        div5            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        div6            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1);
        or3             : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0);
        or4             : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1);
        or5             : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        and3            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1);
        and4            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0);
        and5            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1);
        shl3            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        shl4            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1);
        shl5            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0);
        shr3            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1);
        shr4            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0);
        shr5            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1);
        rol3            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0);
        rol4            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1);
        rol5            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        ror3            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1);
        ror4            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0);
        ror5            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1);
        neg3            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0);
        neg4            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1);
        neg5            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0);
        not3            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi1);
        not4            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0);
        not5            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1);
        ld3             : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0);
        ld4             : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi1);
        ld5             : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0);
        ld6             : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1);
        ld7             : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0);
        ldi3            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1);
        ldi4            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0);
        ldi5            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1);
        st3             : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        st4             : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1);
        st5             : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0);
        st6             : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1);
        st7             : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi0);
        addi3           : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1);
        addi4           : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0);
        addi5           : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1);
        andi3           : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0);
        andi4           : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1);
        andi5           : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0);
        ori3            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1);
        ori4            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0);
        ori5            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        br3             : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        br4             : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        br5             : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        br6             : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1);
        br7             : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        jr3             : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1);
        jal3            : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        jal4            : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1);
        mfhi3           : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        mflo3           : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1);
        in3             : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        out3            : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1);
        nop3            : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0);
        halt3           : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1);
        shra3           : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0);
        shra4           : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1);
        shra5           : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0)
    );
    port(
        HIin            : out    vl_logic;
        LOin            : out    vl_logic;
        PCin            : out    vl_logic;
        MDRin           : out    vl_logic;
        Zin             : out    vl_logic;
        Yin             : out    vl_logic;
        MARin           : out    vl_logic;
        IRin            : out    vl_logic;
        CONin           : out    vl_logic;
        OUTPORTin       : out    vl_logic;
        HIout           : out    vl_logic;
        LOout           : out    vl_logic;
        ZHIout          : out    vl_logic;
        ZLOout          : out    vl_logic;
        PCout           : out    vl_logic;
        MDRout          : out    vl_logic;
        INPORTout       : out    vl_logic;
        OUTPORTout      : out    vl_logic;
        Yout            : out    vl_logic;
        Cout            : out    vl_logic;
        Gra             : out    vl_logic;
        Grb             : out    vl_logic;
        Grc             : out    vl_logic;
        Rin             : out    vl_logic;
        Rout            : out    vl_logic;
        BAout           : out    vl_logic;
        Read            : out    vl_logic;
        IncPC           : out    vl_logic;
        Write           : out    vl_logic;
        Run             : out    vl_logic;
        regIn           : out    vl_logic_vector(15 downto 0);
        Clock           : in     vl_logic;
        Reset           : in     vl_logic;
        Stop            : in     vl_logic;
        IR              : in     vl_logic_vector(31 downto 0);
        present_state   : out    vl_logic_vector(7 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of reset_state : constant is 1;
    attribute mti_svvh_generic_type of fetch0 : constant is 1;
    attribute mti_svvh_generic_type of fetch1 : constant is 1;
    attribute mti_svvh_generic_type of fetch2 : constant is 1;
    attribute mti_svvh_generic_type of add3 : constant is 1;
    attribute mti_svvh_generic_type of add4 : constant is 1;
    attribute mti_svvh_generic_type of add5 : constant is 1;
    attribute mti_svvh_generic_type of sub3 : constant is 1;
    attribute mti_svvh_generic_type of sub4 : constant is 1;
    attribute mti_svvh_generic_type of sub5 : constant is 1;
    attribute mti_svvh_generic_type of mul3 : constant is 1;
    attribute mti_svvh_generic_type of mul4 : constant is 1;
    attribute mti_svvh_generic_type of mul5 : constant is 1;
    attribute mti_svvh_generic_type of mul6 : constant is 1;
    attribute mti_svvh_generic_type of div3 : constant is 1;
    attribute mti_svvh_generic_type of div4 : constant is 1;
    attribute mti_svvh_generic_type of div5 : constant is 1;
    attribute mti_svvh_generic_type of div6 : constant is 1;
    attribute mti_svvh_generic_type of or3 : constant is 1;
    attribute mti_svvh_generic_type of or4 : constant is 1;
    attribute mti_svvh_generic_type of or5 : constant is 1;
    attribute mti_svvh_generic_type of and3 : constant is 1;
    attribute mti_svvh_generic_type of and4 : constant is 1;
    attribute mti_svvh_generic_type of and5 : constant is 1;
    attribute mti_svvh_generic_type of shl3 : constant is 1;
    attribute mti_svvh_generic_type of shl4 : constant is 1;
    attribute mti_svvh_generic_type of shl5 : constant is 1;
    attribute mti_svvh_generic_type of shr3 : constant is 1;
    attribute mti_svvh_generic_type of shr4 : constant is 1;
    attribute mti_svvh_generic_type of shr5 : constant is 1;
    attribute mti_svvh_generic_type of rol3 : constant is 1;
    attribute mti_svvh_generic_type of rol4 : constant is 1;
    attribute mti_svvh_generic_type of rol5 : constant is 1;
    attribute mti_svvh_generic_type of ror3 : constant is 1;
    attribute mti_svvh_generic_type of ror4 : constant is 1;
    attribute mti_svvh_generic_type of ror5 : constant is 1;
    attribute mti_svvh_generic_type of neg3 : constant is 1;
    attribute mti_svvh_generic_type of neg4 : constant is 1;
    attribute mti_svvh_generic_type of neg5 : constant is 1;
    attribute mti_svvh_generic_type of not3 : constant is 1;
    attribute mti_svvh_generic_type of not4 : constant is 1;
    attribute mti_svvh_generic_type of not5 : constant is 1;
    attribute mti_svvh_generic_type of ld3 : constant is 1;
    attribute mti_svvh_generic_type of ld4 : constant is 1;
    attribute mti_svvh_generic_type of ld5 : constant is 1;
    attribute mti_svvh_generic_type of ld6 : constant is 1;
    attribute mti_svvh_generic_type of ld7 : constant is 1;
    attribute mti_svvh_generic_type of ldi3 : constant is 1;
    attribute mti_svvh_generic_type of ldi4 : constant is 1;
    attribute mti_svvh_generic_type of ldi5 : constant is 1;
    attribute mti_svvh_generic_type of st3 : constant is 1;
    attribute mti_svvh_generic_type of st4 : constant is 1;
    attribute mti_svvh_generic_type of st5 : constant is 1;
    attribute mti_svvh_generic_type of st6 : constant is 1;
    attribute mti_svvh_generic_type of st7 : constant is 1;
    attribute mti_svvh_generic_type of addi3 : constant is 1;
    attribute mti_svvh_generic_type of addi4 : constant is 1;
    attribute mti_svvh_generic_type of addi5 : constant is 1;
    attribute mti_svvh_generic_type of andi3 : constant is 1;
    attribute mti_svvh_generic_type of andi4 : constant is 1;
    attribute mti_svvh_generic_type of andi5 : constant is 1;
    attribute mti_svvh_generic_type of ori3 : constant is 1;
    attribute mti_svvh_generic_type of ori4 : constant is 1;
    attribute mti_svvh_generic_type of ori5 : constant is 1;
    attribute mti_svvh_generic_type of br3 : constant is 1;
    attribute mti_svvh_generic_type of br4 : constant is 1;
    attribute mti_svvh_generic_type of br5 : constant is 1;
    attribute mti_svvh_generic_type of br6 : constant is 1;
    attribute mti_svvh_generic_type of br7 : constant is 1;
    attribute mti_svvh_generic_type of jr3 : constant is 1;
    attribute mti_svvh_generic_type of jal3 : constant is 1;
    attribute mti_svvh_generic_type of jal4 : constant is 1;
    attribute mti_svvh_generic_type of mfhi3 : constant is 1;
    attribute mti_svvh_generic_type of mflo3 : constant is 1;
    attribute mti_svvh_generic_type of in3 : constant is 1;
    attribute mti_svvh_generic_type of out3 : constant is 1;
    attribute mti_svvh_generic_type of nop3 : constant is 1;
    attribute mti_svvh_generic_type of halt3 : constant is 1;
    attribute mti_svvh_generic_type of shra3 : constant is 1;
    attribute mti_svvh_generic_type of shra4 : constant is 1;
    attribute mti_svvh_generic_type of shra5 : constant is 1;
end control_unit;

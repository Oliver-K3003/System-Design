/*module multiplier(input signed [31:0] m, input signed [31:0] q, output [63:0] out);

	reg [63:0] product;
	reg [2:0] compare;
	reg []
	
	compare[2] = q[1];
	compare[1] = q[0];
	compare[0] = 1'b0;
	//check the case for the recoding
	case(compare)
		3'b000 : <= //0*M
		3'b001 : <= //+1*M
		3'b010 : <= //+1*M
		3'b011 : <= //+2*M
		3'b100 : <= //-2*M
		3'b101 : <= //-1*M
		3'b110 : <= //-1*M
		3'b111 : <= //0*M
	endcase*/
		
library verilog;
use verilog.vl_types.all;
entity busEncodertb is
end busEncodertb;
